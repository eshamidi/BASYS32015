
Library ieee;
Use ieee.std_logic_1164.all;
Package p1_pack is
Type sh_reg_sel is (no_op, load, shift);
End p1_pack; 